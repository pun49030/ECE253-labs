module part3(Clock, Resetn, Go, Divisor, Dividend, Quotient, Remainder);
	 input Clock;
    input Resetn;
    input Go;
    input [4:0] Divisor;
	 input [3:0] Dividend;
    output [3:0] Quotient;
	 output [4:0] Remainder;
	
module control(
    input clk,
    input resetn,
    input go,

    output reg  ld_a, ld_b, ld_c, ld_x, ld_r,
    output reg  ld_alu_out,
    output reg [1:0]  alu_select_a, alu_select_b,
    output reg alu_op
    );

    reg [5:0] current_state, next_state; 
    

module datapath(
    input clk,
    input resetn,
    input [7:0] data_in,
    input ld_alu_out, 
    input ld_x, ld_a, ld_b, ld_c,
    input ld_r,
    input alu_op, 
    input [1:0] alu_select_a, alu_select_b,
    output reg [7:0] data_result
    );
    